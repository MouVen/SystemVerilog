//https://mouven.blogspot.com/2023/08/wierd-algorithm-in-system-verilog.html

class solution;

    function void your_solution(input bit [63:0] n, ref bit [63:0] q[$]);
      //Type your Solution Here
    endfunction: your_solution

endclass: solution