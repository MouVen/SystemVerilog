//Problem Description: https://mouven.blogspot.com/2023/08/system-verilog-hello-world.html
class solution;

    function void your_solution(output string s);
    //Type your Solution Here
    endfunction

endclass