//Problem Description: <link to blogger>
class solution;
  	function void your_solution(output string s);
    endfunction
endclass